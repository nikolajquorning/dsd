--Tom fil